LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY work;

ENTITY POLARITY_VHDL IS
	PORT
	(
	
		IN_1, IN_2, IN_3, IN_4, POLARITY_CNTRL: IN BIT;
		OUT_1, OUT_2, OUT_3,OUT_4: OUT BIT
		);
END POLARITY_VHDL;

ARCHITECTURE inverter OF POLARITY_VHDL IS

BEGIN

OUT_1 <= IN_1 XOR POLARITY_CNTRL;
OUT_2 <= IN_2 XOR POLARITY_CNTRL;
OUT_3 <= IN_3 XOR POLARITY_CNTRL;
OUT_4 <= IN_4 XOR POLARITY_CNTRL;

END inverter;	
